* SPICE	Mon Apr 29 15:05:39 2024	compleja_def_not
* icv_netlist Version RHEL64 U-2022.12-SP4.9133772 2023/08/28

* Hierarchy Level 0

* Top of hierarchy  cell=compleja_def_not
.subckt compleja_def_not net9 gnd! Out In
X1 Out In gnd! gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.88e-06 ps=1.615e-06
+	 ad=2.064e-13 as=2.3895e-13
X2 gnd! In Out gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.615e-06 ps=1.04e-06
+	 ad=2.3895e-13 as=1.182e-13
X3 Out In gnd! gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.615e-06
+	 ad=1.182e-13 as=2.3895e-13
X4 gnd! In Out gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.615e-06 ps=1.04e-06
+	 ad=2.3895e-13 as=1.182e-13
X5 Out In gnd! gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.615e-06
+	 ad=1.182e-13 as=2.3895e-13
X6 gnd! In Out gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.615e-06 ps=1.04e-06
+	 ad=2.3895e-13 as=1.182e-13
X7 Out In gnd! gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.615e-06
+	 ad=1.182e-13 as=2.3895e-13
X8 gnd! In Out gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.615e-06 ps=1.04e-06
+	 ad=2.3895e-13 as=1.182e-13
X9 Out In gnd! gnd! ne  l=1.8e-07 w=3e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=3.03e-06
+	 ad=1.182e-13 as=4.479e-13
X10 gnd! Out p_dn  area=3.825e-13 pj=2.6e-06 perimeter=2.6e-06
X11 gnd! net9 p_dnw  area=4.85397e-11 pj=3.708e-05 perimeter=3.708e-05
X12 Out In net9 net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.88e-06 ps=1.535e-06
+	 ad=2.164e-13 as=2.3215e-13
X13 net9 In Out net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.535e-06 ps=1.04e-06
+	 ad=2.3215e-13 as=1.282e-13
X14 Out In net9 net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.535e-06
+	 ad=1.282e-13 as=2.3215e-13
X15 net9 In Out net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.535e-06 ps=1.04e-06
+	 ad=2.3215e-13 as=1.282e-13
X16 Out In net9 net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.535e-06
+	 ad=1.282e-13 as=2.3215e-13
X17 net9 In Out net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.535e-06 ps=1.04e-06
+	 ad=2.3215e-13 as=1.282e-13
X18 Out In net9 net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.535e-06
+	 ad=1.282e-13 as=2.3215e-13
X19 net9 In Out net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.535e-06 ps=1.04e-06
+	 ad=2.3215e-13 as=1.282e-13
X20 Out In net9 net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.535e-06
+	 ad=1.282e-13 as=2.3215e-13
X21 net9 In Out net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.535e-06 ps=1.04e-06
+	 ad=2.3215e-13 as=1.282e-13
X22 Out In net9 net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=1.535e-06
+	 ad=1.282e-13 as=2.3215e-13
X23 net9 In Out net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.535e-06 ps=1.04e-06
+	 ad=2.3215e-13 as=1.282e-13
X24 Out In net9 net9 pe  l=1.8e-07 w=4e-07 nrd=-1 nrs=-1 pd=1.04e-06 ps=2.87e-06
+	 ad=1.282e-13 as=4.243e-13
.ends compleja_def_not
